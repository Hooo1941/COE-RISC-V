library verilog;
use verilog.vl_types.all;
entity xgriscv_tb is
end xgriscv_tb;
